library verilog;
use verilog.vl_types.all;
entity top_vlg_tst is
end top_vlg_tst;
